`ifndef DEFINES
`define DEFINES

    //----------------//
    // INSTRN Defines
    //----------------//

    `define INSTRN_CSR(instrn)        (instrn[31:20])
    `define INSTRN_MEM_SIZE(instrn)   (instrn[13:12])
    `define INSTRN_MEM_SIGN(instrn)   (instrn[14])
    `define INSTRN_FM_FENCE(instrn)   (instrn[31:28])

    `define INSTRN_FUNCT7(instrn)     (instrn[31:25])
    `define INSTRN_RS2_ADDR(instrn)   (instrn[24:20])
    `define INSTRN_RS1_ADDR(instrn)   (instrn[19:15])
    `define INSTRN_FUNCT3(instrn)     (instrn[14:12])
    `define INSTRN_RD_ADDR(instrn)    (instrn[11:7])
    `define INSTRN_OPCODE(instrn)     (instrn[6:0])

    // Opcodes
    localparam OPCODE_OP_REG = 7'b0110011;
    localparam OPCODE_OP_IMM = 7'b0010011;
    localparam OPCODE_JALR   = 7'b1100111;
    localparam OPCODE_LOAD   = 7'b0000011;
    localparam OPCODE_STORE  = 7'b0100011;
    localparam OPCODE_BRANCH = 7'b1100011;
    localparam OPCODE_LUI    = 7'b0110111;
    localparam OPCODE_AUIPC  = 7'b0010111;
    localparam OPCODE_JAL    = 7'b1101111;
    localparam OPCODE_FENCE  = 7'b0001111;
    localparam OPCODE_SYS    = 7'b1110011;

    // Opcode FUNCT3s
    localparam FUNCT3_I_JALR    = 3'b000;

    localparam FUNCT3_I_LB      = 3'b000;
    localparam FUNCT3_I_LH      = 3'b001;
    localparam FUNCT3_I_LW      = 3'b010;
    localparam FUNCT3_I_LBU     = 3'b100;
    localparam FUNCT3_I_LHU     = 3'b101;

    localparam FUNCT3_I_ADDI    = 3'b000;
    localparam FUNCT3_I_SLTI    = 3'b010;
    localparam FUNCT3_I_SLTIU   = 3'b011;
    localparam FUNCT3_I_ORI     = 3'b110;
    localparam FUNCT3_I_XORI    = 3'b100;
    localparam FUNCT3_I_ANDI    = 3'b111;
    localparam FUNCT3_I_SLI     = 3'b001;
    localparam FUNCT3_I_SRI     = 3'b101;

    localparam FUNCT3_B_BEQ     = 3'b000;
    localparam FUNCT3_B_BNE     = 3'b001;
    localparam FUNCT3_B_BLT     = 3'b100;
    localparam FUNCT3_B_BGE     = 3'b101;
    localparam FUNCT3_B_BLTU    = 3'b110;
    localparam FUNCT3_B_BGEU    = 3'b111;

    localparam FUNCT3_S_SB      = 3'b000;
    localparam FUNCT3_S_SH      = 3'b001;
    localparam FUNCT3_S_SW      = 3'b010;

    localparam FUNCT3_R_ADD     = 3'b000;
    localparam FUNCT3_R_SUB     = 3'b000;
    localparam FUNCT3_R_SLL     = 3'b001;
    localparam FUNCT3_R_SLT     = 3'b010;
    localparam FUNCT3_R_SLTU    = 3'b011;
    localparam FUNCT3_R_XOR     = 3'b100;
    localparam FUNCT3_R_SRL     = 3'b101;
    localparam FUNCT3_R_SRA     = 3'b101;
    localparam FUNCT3_R_OR      = 3'b110;
    localparam FUNCT3_R_AND     = 3'b111;

    localparam FUNCT3_FENCE     = 3'b000;
    localparam FUNCT3_FENCE_I   = 3'b001;

    localparam FUNCT3_SYS_CSRRW  = 3'b001;
    localparam FUNCT3_SYS_CSRRS  = 3'b010;
    localparam FUNCT3_SYS_CSRRC  = 3'b011;
    localparam FUNCT3_SYS_CSRRWI = 3'b101;
    localparam FUNCT3_SYS_CSRRSI = 3'b110;
    localparam FUNCT3_SYS_CSRRCI = 3'b111;
    localparam FUNCT3_SYS_TRAPS  = 3'b000;

    // Instruction FUNCT7s
    localparam FUNCT7_I_R_Z = 7'bzzzzzzz;
    localparam FUNCT7_I_R_0 = 7'b0000000;
    localparam FUNCT7_I_R_1 = 7'b0100000;

    localparam FUNCT7_RS2_SYS_ECALL  = 12'h000;
    localparam FUNCT7_RS2_SYS_EBREAK = 12'h001;
    localparam FUNCT7_RS2_SYS_MRET   = 12'h302;
    localparam FUNCT7_RS2_SYS_WFI    = 12'h205;

    localparam FM_FENCE              = 4'bz000;

    //--------------//
    // ALU Defines
    //--------------//

    localparam ALU_ADD  = 4'b0000;
    localparam ALU_SUB  = 4'b1000;
    localparam ALU_OR   = 4'b0110;
    localparam ALU_AND  = 4'b0111;
    localparam ALU_XOR  = 4'b0100;
    localparam ALU_SRL  = 4'b0101;
    localparam ALU_SLL  = 4'b0001;
    localparam ALU_SRA  = 4'b1101;
    localparam ALU_SLT  = 4'b0010;
    localparam ALU_SLTU = 4'b0011;
    localparam ALU_LUI  = 4'b1001;

    localparam ALU_SRC_SEL_A_RS1       = 1'd0;
    localparam ALU_SRC_SEL_A_UPPER_IMM = 1'd1;

    localparam ALU_SRC_SEL_B_RS2         = 2'd0;
    localparam ALU_SRC_SEL_B_I_TYPE_IMM  = 2'd1;
    localparam ALU_SRC_SEL_B_S_TYPE_IMM  = 2'd2;
    localparam ALU_SRC_SEL_B_PC_ADDR     = 2'd3;

    //--------------//
    // CSR Defines
    //--------------//

    // Read-Only Addresses
    localparam CSR_MVENDORID_ADDR  = 12'hF11;
    localparam CSR_MARCHID_ADDR    = 12'hF12;
    localparam CSR_MIMPID_ADDR     = 12'hF13;
    localparam CSR_MHARTID_ADDR    = 12'hF14;
    localparam CSR_MCONFIGPTR_ADDR = 12'hF15;

    // Trap Addresses
    localparam CSR_MSTATUS_ADDR  = 12'h300;
    localparam CSR_MISA_ADDR     = 12'h301;
    localparam CSR_MIE_ADDR      = 12'h304;
    localparam CSR_MTVEC_ADDR    = 12'h305;
    localparam CSR_MSTATUSH_ADDR = 12'h310;
    localparam CSR_MSCRATCH_ADDR = 12'h340;
    localparam CSR_MEPC_ADDR     = 12'h341;
    localparam CSR_MCAUSE_ADDR   = 12'h342;
    localparam CSR_MTVAL_ADDR    = 12'h343;
    localparam CSR_MIP_ADDR      = 12'h344;


	localparam CSR_MCYCLE_ADDR    = 12'hB00;
	localparam CSR_MINSTRET_ADDR  = 12'hB02;
	localparam CSR_MCYCLEH_ADDR   = 12'hB80;
	localparam CSR_MINSTRETH_ADDR = 12'hB82;


    // MCAUSE Codes
    localparam MCAUSE_SEL_NOP                  = 3'd0;
    localparam MCAUSE_SEL_INSTRN_ADDR_MISALIGN = 3'd1;
    localparam MCAUSE_SEL_INVLD_INSTRN         = 3'd2;
    localparam MCAUSE_SEL_LOAD_ADDR_MISALIGN   = 3'd3;
    localparam MCAUSE_SEL_STORE_ADDR_MISALIGN  = 3'd4;

    localparam MCAUSE_CODE_INSTRN_ADDR_MISALIGN = 32'h00000000;
    localparam MCAUSE_CODE_INVLD_INSTRN         = 32'h00000002;
    localparam MCAUSE_CODE_BREAKPOINT           = 32'h00000003;
    localparam MCAUSE_CODE_LOAD_ADDR_MISALIGN   = 32'h00000004;
    localparam MCAUSE_CODE_STORE_ADDR_MISALIGN  = 32'h00000006;
    localparam MCAUSE_CODE_ECALL_M_MODE         = 32'h0000000b;

    localparam MCAUSE_CODE_MACHINE_SOFTWARE_INTERRUPT = 32'h80000003;
    localparam MCAUSE_CODE_MACHINE_TIMER_INTERRUPT    = 32'h80000007;
    localparam MCAUSE_CODE_MACHINE_EXTERNAL_INTERRUPT = 32'h8000000b;

    // CSR Func Selectors
    localparam CSR_OP_WRITE  = 3'd0;
    localparam CSR_OP_ECALL  = 3'd1;
    localparam CSR_OP_EBREAK = 3'd2;
    localparam CSR_OP_MRET   = 3'd3;
    localparam CSR_OP_WFI    = 3'd4;
    localparam CSR_OP_INTRPT = 3'd5;
    localparam CSR_OP_TRAP   = 3'd6;
    localparam CSR_OP_RESET  = 3'd7;

    localparam CSR_FUNCT3_LOW_RW = 2'b01;
    localparam CSR_FUNCT3_LOW_RS = 2'b10;
    localparam CSR_FUNCT3_LOW_RC = 2'b11;
    localparam CSR_FUNCT3_HIGH_REG = 1'b0;
    localparam CSR_FUNCT3_HIGH_IMM = 1'b1;

    //--------------//
    // MEM Defines
    //--------------//

    localparam MEM_SIZE_BYTE   = 2'd0;
    localparam MEM_SIZE_H_WORD = 2'd1;
    localparam MEM_SIZE_WORD   = 2'd2;

    //--------------//
    // RFILE Defines
    //--------------//

    localparam RFILE_W_SEL_PC_ADDR_INC  = 2'd0;
    localparam RFILE_W_SEL_CSR_R_DATA   = 2'd1;
    localparam RFILE_W_SEL_DMEM_R_DATA  = 2'd2;
    localparam RFILE_W_SEL_ALU_RESULT   = 2'd3;

    //--------------//
    // PC Defines
    //--------------//

    localparam PC_SRC_SEL_ADDR_INC  = 3'd0;
    localparam PC_SRC_SEL_JALR      = 3'd1;
    localparam PC_SRC_SEL_BRANCH    = 3'd2;
    localparam PC_SRC_SEL_JAL       = 3'd3;
    localparam PC_SRC_SEL_MTVEC     = 3'd4;
    localparam PC_SRC_SEL_MEPC      = 3'd5;
    localparam PC_SRC_SEL_RESET_VEC = 3'd6;

    //--------------//
    // FSM Defines
    //--------------//

    localparam ST_INIT   = 2'd0;
    localparam ST_EXEC   = 2'd1;
    localparam ST_WR_BK  = 2'd2;

    //--------------//
    // RVFI Defines
    //--------------//

    `define RVFI_CSR_LIST \
        `CSR_MACRO_OP(mstatus)    \
        `CSR_MACRO_OP(misa)       \
        `CSR_MACRO_OP(mie)        \
        `CSR_MACRO_OP(mtvec)      \
        `CSR_MACRO_OP(mstatush)   \
        `CSR_MACRO_OP(mscratch)   \
        `CSR_MACRO_OP(mepc)       \
        `CSR_MACRO_OP(mcause)     \
        `CSR_MACRO_OP(mtval)      \
        `CSR_MACRO_OP(mip)        \
        `CSR_MACRO_OP(mvendorid)  \
        `CSR_MACRO_OP(marchid)    \
        `CSR_MACRO_OP(mimpid)     \
        `CSR_MACRO_OP(mhartid)    \
        `CSR_MACRO_OP(mconfigptr)

    `define CSR_MACRO_OP(NAME) \
        output reg [31:0] rvfi_csr_``NAME``_rmask, \
        output reg [31:0] rvfi_csr_``NAME``_wmask, \
        output reg [31:0] rvfi_csr_``NAME``_rdata, \
        output reg [31:0] rvfi_csr_``NAME``_wdata,
    `undef CSR_MACRO_OP

    // Assignments
    `define CSR_MACRO_OP(NAME) \
        rvfi_csr_``NAME``_rmask <= 32'hffff_ffff; \
        rvfi_csr_``NAME``_wmask <= 32'hffff_ffff; \
        rvfi_csr_``NAME``_rdata <= csr_``NAME``; \
        rvfi_csr_``NAME``_wdata <= csr_``NAME``;
    `undef CSR_MACRO_OP

    `define RVFI_OUTPUTS                  \
        output reg        rvfi_valid,     \
        output reg [63:0] rvfi_order,     \
        output reg [31:0] rvfi_insn,      \
        output reg        rvfi_trap,      \
        output reg        rvfi_halt,      \
        output reg        rvfi_intr,      \
        output reg [ 1:0] rvfi_mode,      \
        output reg [ 1:0] rvfi_ixl,       \
        output reg [ 4:0] rvfi_rs1_addr,  \
        output reg [ 4:0] rvfi_rs2_addr,  \
        output reg [31:0] rvfi_rs1_rdata, \
        output reg [31:0] rvfi_rs2_rdata, \
        output reg [ 4:0] rvfi_rd_addr,   \
        output reg [31:0] rvfi_rd_wdata,  \
        output reg [31:0] rvfi_pc_rdata,  \
        output reg [31:0] rvfi_pc_wdata,  \
        output reg [31:0] rvfi_mem_addr,  \
        output reg [ 3:0] rvfi_mem_rmask, \
        output reg [ 3:0] rvfi_mem_wmask, \
        output reg [31:0] rvfi_mem_rdata, \
        output reg [31:0] rvfi_mem_wdata, \
        `RVFI_CSR_LIST

`endif
