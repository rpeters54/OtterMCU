`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/02/2022 03:54:39 PM
// Desmode 
// Module Name: CU_DCDR
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`include "otter_defines.vh"

module otter_cu_dcdr (
    input            clk,
    input            rst,
    input     [31:0] instrn,

    // Branch Signals
    input            br_eq, 
    input            br_lt, 
    input            br_ltu,

    // CSR Signals
    input            csr_intrpt_vld,
    input            csr_addr_vld,
    input            csr_read_only,

    // Alignment Signals
    input      [1:0] addr_store_alignment,
    input      [1:0] addr_load_alignment,
    input      [1:0] addr_jalr_alignment,
    input      [1:0] addr_branch_alignment,
    input      [1:0] addr_jal_alignment,

    // stateless outputs (dependent on decoded inst)
    output reg [3:0] alu_func,
    output reg       alu_src_sel_a,
    output reg [1:0] alu_src_sel_b,
    output reg [1:0] rfile_w_sel,
    output reg [2:0] pc_src_sel,
    output reg [2:0] csr_op_sel,
    output reg [3:0] dmem_w_strb,

    // stateful outputs (dependent on fsm)
    output reg        pc_w_en, 
    output reg        rfile_w_en,
    output reg        dmem_w_en,
    output reg        dmem_r_en,
    output reg        csr_w_en,
    output reg        stall
);

    reg illegal_instrn, write_attempt;

    // decompose instruction into component parts
    wire [6:0] funct7   = `INSTRN_FUNCT7(instrn);
    wire [4:0] rs2_addr = `INSTRN_RS2_ADDR(instrn);
    wire [4:0] rs1_addr = `INSTRN_RS1_ADDR(instrn);
    wire [2:0] funct3   = `INSTRN_FUNCT3(instrn);
    wire [4:0] rd_addr  = `INSTRN_RD_ADDR(instrn);
    wire [6:0] opcode   = `INSTRN_OPCODE(instrn);

    // state variables and initial values
    reg [2:0] present_state, next_state;
    initial begin
        present_state = ST_INIT;
	    next_state    = ST_INIT;
    end

    // state update block
    always @(posedge clk) begin
        if (rst == '1) begin
            present_state <= ST_INIT;
        end else begin
            present_state <= next_state;
        end
    end


    always @(*) begin

        // stateless defaults
        alu_func        = ALU_ADD; 
        alu_src_sel_a   = ALU_SRC_SEL_A_RS1; 
        alu_src_sel_b   = ALU_SRC_SEL_B_RS2;
        rfile_w_sel     = RFILE_W_SEL_PC_ADDR_INC; 
        pc_src_sel      = PC_SRC_SEL_ADDR_INC; 
        csr_op_sel      = CSR_OP_WRITE;
        illegal_instrn  = '0;

        // stateful defaults
        pc_w_en      = '1; 
        rfile_w_en   = '0; 
        dmem_w_en    = '0; 
        dmem_r_en    = '0; 
        csr_w_en     = '0; 
        stall        = '0;

        case (present_state)
            ST_INIT : begin
                pc_w_en    = '0; 
                stall      = '1; 
                next_state = ST_EXEC;
            end
            ST_EXEC :  begin
                next_state = ST_EXEC;

                case(opcode)
                    OPCODE_OP_REG : begin    // R-Type opcode
                        case ({funct7, funct3})  // arithmetic/logical operations including two registers
                            {FUNCT7_I_R_0, FUNCT3_R_ADD},
                            {FUNCT7_I_R_1, FUNCT3_R_SUB}, 
                            {FUNCT7_I_R_0, FUNCT3_R_SLL},
                            {FUNCT7_I_R_0, FUNCT3_R_SLT},
                            {FUNCT7_I_R_0, FUNCT3_R_SLTU},
                            {FUNCT7_I_R_0, FUNCT3_R_XOR},
                            {FUNCT7_I_R_0, FUNCT3_R_SRL},
                            {FUNCT7_I_R_1, FUNCT3_R_SRA},
                            {FUNCT7_I_R_0, FUNCT3_R_OR},
                            {FUNCT7_I_R_0, FUNCT3_R_AND} : begin
                                alu_src_sel_a = ALU_SRC_SEL_A_RS1;
                                alu_src_sel_b = ALU_SRC_SEL_B_RS2;
                                rfile_w_sel   = RFILE_W_SEL_ALU_RESULT;
                                alu_func      = {instrn[30], funct3}; 

                                rfile_w_en = '1;
                            end
                            default begin 
                                illegal_instrn = '1;
                            end
                        endcase
                    end
                    OPCODE_OP_IMM : begin    // I-Type opcode *no loading
                        casez ({funct7, funct3}) // arithmetic/logical operations including a register and immediate
                            {FUNCT7_I_R_Z, FUNCT3_I_ADDI},
                            {FUNCT7_I_R_Z, FUNCT3_I_SLTI}, 
                            {FUNCT7_I_R_Z, FUNCT3_I_SLTIU}, 
                            {FUNCT7_I_R_Z, FUNCT3_I_ORI},
                            {FUNCT7_I_R_Z, FUNCT3_I_XORI}, 
                            {FUNCT7_I_R_Z, FUNCT3_I_ANDI}, 
                            {FUNCT7_I_R_0, FUNCT3_I_SLI}, 
                            {FUNCT7_I_R_0, FUNCT3_I_SRI},
                            {FUNCT7_I_R_1, FUNCT3_I_SRI} : begin
                                alu_src_sel_a = ALU_SRC_SEL_A_RS1; 
                                alu_src_sel_b = ALU_SRC_SEL_B_I_TYPE_IMM;
                                rfile_w_sel   = RFILE_W_SEL_ALU_RESULT;
                                alu_func      = {(funct3 == FUNCT3_I_SRI) && instrn[30], funct3};

                                rfile_w_en = '1;
                            end
                            default begin 
                                illegal_instrn = '1;
                            end
                        endcase
                    end
                    OPCODE_JALR : begin    // I-Type opcode *jalr
                        if (funct3 == FUNCT3_I_JALR && addr_jalr_alignment == 2'b00) begin
                            rfile_w_sel = RFILE_W_SEL_PC_ADDR_INC;
                            pc_src_sel  = PC_SRC_SEL_JALR;

                            rfile_w_en = '1;
                        end else begin
                            illegal_instrn = '1;
                        end
                    end
                    OPCODE_LOAD : begin      // I-Type opcode *load instructions
                        alu_src_sel_a = ALU_SRC_SEL_A_RS1;
                        alu_src_sel_b = ALU_SRC_SEL_B_I_TYPE_IMM;
                        alu_func      = ALU_ADD;

                        // Note: alu_result is the computed address
                        casez ({funct3, addr_load_alignment})
                            {FUNCT3_I_LB,  2'bzz},
                            {FUNCT3_I_LH,  2'bz0}, 
                            {FUNCT3_I_LW,  2'b00},
                            {FUNCT3_I_LBU, 2'bzz}, 
                            {FUNCT3_I_LHU, 2'bz0} : begin

                                dmem_r_en  = '1;
                                pc_w_en    = '0;
                                stall      = '1; 
                                next_state = ST_WR_BK;
                            end
                            default begin 
                                illegal_instrn = '1;
                            end
                        endcase
                    end
                    OPCODE_STORE : begin     // S-Type opcode *store instructions
                        alu_src_sel_a = ALU_SRC_SEL_A_RS1; 
                        alu_src_sel_b = ALU_SRC_SEL_B_S_TYPE_IMM;
                        alu_func      = ALU_ADD;

                        // Note: alu_result is the computed address
                        casez ({funct3, addr_store_alignment})
                            {FUNCT3_S_SB, 2'bzz},
                            {FUNCT3_S_SH, 2'bz0},
                            {FUNCT3_S_SW, 2'b00} : begin

                                dmem_w_strb = 4'b 1111;
                                case (funct3)
                                    FUNCT3_S_SB : dmem_w_strb = 4'b 0001;
                                    FUNCT3_S_SH : dmem_w_strb = 4'b 0011;
                                    FUNCT3_S_SW : dmem_w_strb = 4'b 1111;
                                    default : ;
                                endcase
                                // shift to handle different byte/nibble alignments
                                dmem_w_strb = dmem_w_strb << addr_store_alignment;

                                dmem_w_en = '1;
                            end
                            default begin 
                                illegal_instrn = '1;
                            end
                        endcase
                    end
                    OPCODE_BRANCH : begin  // B-Type opcode
                        case (funct3) // All store instructions; writing from registers to memory
                            FUNCT3_B_BEQ, FUNCT3_B_BNE, FUNCT3_B_BLT,
                            FUNCT3_B_BGE, FUNCT3_B_BLTU, FUNCT3_B_BGEU : begin
                                if ( // branch taken
                                    (funct3 == FUNCT3_B_BEQ  &&  br_eq)  ||
                                    (funct3 == FUNCT3_B_BNE  && !br_eq)  ||
                                    (funct3 == FUNCT3_B_BLT  &&  br_lt)  ||
                                    (funct3 == FUNCT3_B_BGE  && !br_lt)  ||
                                    (funct3 == FUNCT3_B_BLTU &&  br_ltu) ||
                                    (funct3 == FUNCT3_B_BGEU && !br_ltu)
                                ) begin
                                    // only mark misaligned address if branch
                                    // taken (as per spec)
                                    if (addr_branch_alignment  == 2'b00) begin
                                        pc_src_sel = PC_SRC_SEL_BRANCH;
                                    end else begin
                                        illegal_instrn = '1;
                                    end
                                end
                            end
                            default begin
                                illegal_instrn = '1;
                            end
                        endcase
                    end
                    OPCODE_LUI : begin
                        alu_src_sel_a = ALU_SRC_SEL_A_UPPER_IMM; // Extends a 20-bit immediate (extra 12-bits after)
                        rfile_w_sel   = RFILE_W_SEL_ALU_RESULT;
                        alu_func      = ALU_LUI;                     // Value passes through ALU and is stored in a register

                        rfile_w_en = '1;
                    end
                    OPCODE_AUIPC : begin
                        alu_src_sel_a = ALU_SRC_SEL_A_UPPER_IMM; // Adds a U-type immediate to the program count
                        alu_src_sel_b = ALU_SRC_SEL_B_PC_ADDR;   // which is stored in a register
                        rfile_w_sel   = RFILE_W_SEL_ALU_RESULT;
                        alu_func      = ALU_ADD;

                        rfile_w_en = '1;
                    end
                    OPCODE_JAL : begin
                        if (addr_jal_alignment == 2'b00) begin
                            rfile_w_sel = RFILE_W_SEL_PC_ADDR_INC; // stores current location + 4 in a register
                            pc_src_sel  = PC_SRC_SEL_JAL;          // Jumps to a new location (updates PC value)

                            rfile_w_en = '1;
                        end else begin
                            illegal_instrn = '1;
                        end
                    end
                    OPCODE_FENCE : begin
                        casez ({funct7, rs2_addr, rs1_addr, funct3, rd_addr})
                            PREFIX_FENCE, PREFIX_FENCE_I : begin
                                // nop
                            end
                            default : begin
                                illegal_instrn = '1;
                            end
                        endcase
                    end
                    OPCODE_SYS : begin
                        case (funct3)
                            FUNCT3_SYS_CSRRW, FUNCT3_SYS_CSRRS, FUNCT3_SYS_CSRRC, 
                            FUNCT3_SYS_CSRRWI, FUNCT3_SYS_CSRRSI, FUNCT3_SYS_CSRRCI : begin

                                // Values shared between all CSR instructions
                                rfile_w_sel = RFILE_W_SEL_CSR_R_DATA;
                                rfile_w_en = '1;

                                // CSRRS and CSRRC are read-only compatible if rs1 is x0
                                write_attempt = (funct3 == FUNCT3_SYS_CSRRW)
                                    || (funct3 == FUNCT3_SYS_CSRRWI) 
                                    || (rs1_addr != 5'b0);

                                // illegal if csr dne or write to read-only
                                if (!csr_addr_vld || (write_attempt && csr_read_only)) begin
                                    illegal_instrn = 1'b1;
                                end else begin
                                    rfile_w_sel = RFILE_W_SEL_CSR_R_DATA;
                                    rfile_w_en  = 1'b1;
                                    csr_w_en    = write_attempt;
                                    csr_op_sel  = CSR_OP_WRITE;
                                end
                            end
                            FUNCT3_SYS_TRAPS : begin
                                case ({funct7, rs2_addr})
                                    FUNCT7_RS2_SYS_ECALL : begin
                                        pc_src_sel = PC_SRC_SEL_MTVEC;
                                        csr_op_sel = CSR_OP_ECALL;
                                    end
                                    FUNCT7_RS2_SYS_EBREAK : begin
                                        pc_src_sel = PC_SRC_SEL_MTVEC;
                                        csr_op_sel = CSR_OP_EBREAK;
                                    end
                                    FUNCT7_RS2_SYS_MRET : begin
                                        pc_src_sel = PC_SRC_SEL_MEPC;
                                        csr_op_sel = CSR_OP_MRET;
                                    end
                                    FUNCT7_RS2_SYS_WFI : begin
                                        // TODO: make this more than just
                                        // a nop
                                        csr_op_sel = CSR_OP_WFI;
                                    end
                                    default begin
                                        illegal_instrn = '1;
                                    end
                                endcase
                            end
                            default : begin 
                                illegal_instrn = '1;
                            end
                        endcase
                    end
                    default : begin 
                        illegal_instrn = '1;
                    end
                endcase

                // trap case
                if (illegal_instrn) begin
                    pc_src_sel = PC_SRC_SEL_MTVEC;
                    csr_op_sel = CSR_OP_TRAP;
                // interrupt case
                end else if (csr_intrpt_vld) begin
                    pc_src_sel = PC_SRC_SEL_MTVEC;
                    csr_op_sel = CSR_OP_INTRPT;
                end 

                // Avoid writing back if interrupt/trap occurs
                if (csr_intrpt_vld || illegal_instrn) begin
                    pc_w_en      = '1; 
                    rfile_w_en   = '0; 
                    dmem_w_en    = '0; 
                    dmem_r_en    = '0; 
                    csr_w_en     = '0; 
                    stall        = '0; 

                    next_state = ST_EXEC;
                end
            end
            ST_WR_BK : begin
                // memory reads require an extra clock cycle
                rfile_w_sel = RFILE_W_SEL_DMEM_R_DATA;
                rfile_w_en  = '1;
                next_state  = ST_EXEC;
            end
            default : begin 
                next_state = ST_INIT;
            end
        endcase
    end


`ifdef FORMAL

    // Helper signals for formal properties
    wire f_exception_taken = illegal_instrn || csr_intrpt_vld;
    reg  f_past_valid;
    reg  f_past_rst;
    reg [31:0] f_prev_instrn;

    initial begin
        f_past_valid = 0;
        f_past_rst = 0;
        f_prev_cycle_was_load = 0;
        f_prev_instrn = '0;
    end

    always @(posedge clk) begin
        f_past_valid <= 1;
        f_past_rst   <= rst;
        f_prev_instrn <= instrn;
    end

    // --- Assumptions ---
    always @(*) begin
        if (!f_past_valid) assume(rst);
    end

    // --- Assertions ---
    always @(*) begin
        // Property: On reset, the FSM must be in the INIT state.
        if (f_past_rst) assert(present_state == ST_INIT);

        // Property: A trap must take priority over an interrupt.
        if (present_state == ST_EXEC && illegal_instrn)
            assert(csr_op_sel != CSR_OP_INTRPT);

        // Property: When any trap or interrupt is taken, architectural state writes must be disabled.
        if (present_state == ST_EXEC && f_exception_taken)
            assert(pc_w_en       == '1 &&
                   rfile_w_en    == '0 &&
                   dmem_w_en     == '0 &&
                   dmem_r_en     == '0 &&
                   csr_w_en      == '0 &&
                   stall         == '0);

        // R-Type Control Signals
        if (present_state == ST_EXEC && opcode == OPCODE_OP_REG && !f_exception_taken)
            assert(alu_src_sel_a == ALU_SRC_SEL_A_RS1 &&
                   alu_src_sel_b == ALU_SRC_SEL_B_RS2 &&
                   rfile_w_sel   == RFILE_W_SEL_ALU_RESULT &&
                   alu_func      == {instrn[30], funct3} &&
                   pc_src_sel    == PC_SRC_SEL_ADDR_INC &&
                   pc_w_en       == '1 &&
                   rfile_w_en    == '1 &&
                   dmem_w_en     == '0 &&
                   dmem_r_en     == '0 &&
                   csr_w_en      == '0 &&
                   stall         == '0);

        // I-Type Control Signals
        if (present_state == ST_EXEC && opcode == OPCODE_OP_IMM && !f_exception_taken)
            assert(alu_src_sel_a == ALU_SRC_SEL_A_RS1 &&
                   alu_src_sel_b == ALU_SRC_SEL_B_I_TYPE_IMM &&
                   rfile_w_sel   == RFILE_W_SEL_ALU_RESULT &&
                   alu_func      == {(funct3 == FUNCT3_I_SRI) && instrn[30], funct3} &&
                   pc_src_sel    == PC_SRC_SEL_ADDR_INC &&
                   pc_w_en       == '1 &&
                   rfile_w_en    == '1 &&
                   dmem_w_en     == '0 &&
                   dmem_r_en     == '0 &&
                   csr_w_en      == '0 &&
                   stall         == '0);

        // JALR Control Signals
        if (present_state == ST_EXEC && opcode == OPCODE_JALR && !f_exception_taken)
            assert(rfile_w_sel   == RFILE_W_SEL_PC_ADDR_INC &&
                   pc_src_sel    == PC_SRC_SEL_JALR &&
                   pc_w_en       == '1 &&
                   rfile_w_en    == '1 &&
                   dmem_w_en     == '0 &&
                   dmem_r_en     == '0 &&
                   csr_w_en      == '0 &&
                   stall         == '0);

        // Property: For any valid LOAD instruction (first cycle).
        if (present_state == ST_EXEC && opcode == OPCODE_LOAD && !f_exception_taken)
            assert(next_state == ST_WR_BK &&
                   pc_w_en       == '0 &&
                   rfile_w_en    == '0 &&
                   dmem_w_en     == '0 &&
                   dmem_r_en     == '1 &&
                   csr_w_en      == '0 &&
                   stall         == '1);

        if (present_state == ST_WR_BK)
            assert(next_state    == ST_EXEC &&
                   pc_w_en       == '1 &&
                   rfile_w_en    == '1 &&
                   dmem_w_en     == '0 &&
                   dmem_r_en     == '0 &&
                   csr_w_en      == '0 &&
                   stall         == '0);

        // Property: For any valid STORE instruction.
        if (present_state == ST_EXEC && opcode == OPCODE_STORE && !f_exception_taken)
            assert(pc_w_en       == '1 &&
                   rfile_w_en    == '0 &&
                   dmem_w_en     == '1 &&
                   dmem_r_en     == '0 &&
                   csr_w_en      == '0 &&
                   stall         == '0);

        // Property: For a JAL instruction.
        if (present_state == ST_EXEC && opcode == OPCODE_JAL && !f_exception_taken)
            assert(pc_src_sel == PC_SRC_SEL_JAL && rfile_w_en == 1'b1 && rfile_w_sel == RFILE_W_SEL_PC_ADDR_INC);

        // Property: For an ECALL instruction.
        if (present_state == ST_EXEC && instrn == 32'h00000073 && !f_exception_taken) // Full ECALL encoding
            assert(csr_op_sel == CSR_OP_ECALL && pc_src_sel == PC_SRC_SEL_MTVEC);
    end

    // --- Coverage Checks ---
    always @(posedge clk) begin
        cover(present_state == ST_EXEC && opcode == OPCODE_OP_REG && !f_exception_taken);
        cover(present_state == ST_EXEC && opcode == OPCODE_LOAD && !f_exception_taken);
        cover(present_state == ST_EXEC && opcode == OPCODE_STORE && !f_exception_taken);
        cover(present_state == ST_EXEC && opcode == OPCODE_JAL && !f_exception_taken);
        cover(present_state == ST_EXEC && illegal_instrn);
        cover(present_state == ST_EXEC && !illegal_instrn && csr_intrpt_vld);
    end
`endif

endmodule
